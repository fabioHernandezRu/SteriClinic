// mi_nios.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module mi_nios (
		output wire        bl_n_export,       //       bl_n.export
		output wire        bl_p_export,       //       bl_p.export
		input  wire        clk_clk,           //        clk.clk
		output wire        flash_dclk,        //      flash.dclk
		output wire        flash_sce,         //           .sce
		output wire        flash_sdo,         //           .sdo
		input  wire        flash_data0,       //           .data0
		inout  wire [15:0] lcd32_data_export, // lcd32_data.export
		output wire        lcd_cs_export,     //     lcd_cs.export
		output wire        lcd_rd_export,     //     lcd_rd.export
		output wire        lcd_rs_export,     //     lcd_rs.export
		output wire        lcd_wr_export,     //     lcd_wr.export
		output wire [7:0]  led_export,        //        led.export
		input  wire        reset_reset_n,     //      reset.reset_n
		output wire        reset_1_export,    //    reset_1.export
		output wire [11:0] sdram_addr,        //      sdram.addr
		output wire [1:0]  sdram_ba,          //           .ba
		output wire        sdram_cas_n,       //           .cas_n
		output wire        sdram_cke,         //           .cke
		output wire        sdram_cs_n,        //           .cs_n
		inout  wire [15:0] sdram_dq,          //           .dq
		output wire [1:0]  sdram_dqm,         //           .dqm
		output wire        sdram_ras_n,       //           .ras_n
		output wire        sdram_we_n,        //           .we_n
		output wire        sdram_clk_clk,     //  sdram_clk.clk
		input  wire        spi_touch_MISO,    //  spi_touch.MISO
		output wire        spi_touch_MOSI,    //           .MOSI
		output wire        spi_touch_SCLK,    //           .SCLK
		output wire        spi_touch_SS_n,    //           .SS_n
		input  wire [3:0]  sw_export,         //         sw.export
		output wire        touch_cs_export,   //   touch_cs.export
		input  wire        touch_irq_export   //  touch_irq.export
	);

	wire         pll_c0_clk;                                              // pll:c0 -> [bl_n:clk, bl_p:clk, flash:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, lcd32_data:clk, lcd_cs:clk, lcd_rd:clk, lcd_rs:clk, lcd_wr:clk, mm_interconnect_0:pll_c0_clk, niosGe:clk, reset:clk, rst_controller_001:clk, rst_controller_002:clk, sdram:clk, spi_touch:clk, sysid:clock, touch_cs:clk, touch_irq:clk]
	wire  [31:0] niosge_data_master_readdata;                             // mm_interconnect_0:niosGe_data_master_readdata -> niosGe:d_readdata
	wire         niosge_data_master_waitrequest;                          // mm_interconnect_0:niosGe_data_master_waitrequest -> niosGe:d_waitrequest
	wire         niosge_data_master_debugaccess;                          // niosGe:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:niosGe_data_master_debugaccess
	wire  [24:0] niosge_data_master_address;                              // niosGe:d_address -> mm_interconnect_0:niosGe_data_master_address
	wire   [3:0] niosge_data_master_byteenable;                           // niosGe:d_byteenable -> mm_interconnect_0:niosGe_data_master_byteenable
	wire         niosge_data_master_read;                                 // niosGe:d_read -> mm_interconnect_0:niosGe_data_master_read
	wire         niosge_data_master_readdatavalid;                        // mm_interconnect_0:niosGe_data_master_readdatavalid -> niosGe:d_readdatavalid
	wire         niosge_data_master_write;                                // niosGe:d_write -> mm_interconnect_0:niosGe_data_master_write
	wire  [31:0] niosge_data_master_writedata;                            // niosGe:d_writedata -> mm_interconnect_0:niosGe_data_master_writedata
	wire  [31:0] niosge_instruction_master_readdata;                      // mm_interconnect_0:niosGe_instruction_master_readdata -> niosGe:i_readdata
	wire         niosge_instruction_master_waitrequest;                   // mm_interconnect_0:niosGe_instruction_master_waitrequest -> niosGe:i_waitrequest
	wire  [24:0] niosge_instruction_master_address;                       // niosGe:i_address -> mm_interconnect_0:niosGe_instruction_master_address
	wire         niosge_instruction_master_read;                          // niosGe:i_read -> mm_interconnect_0:niosGe_instruction_master_read
	wire         niosge_instruction_master_readdatavalid;                 // mm_interconnect_0:niosGe_instruction_master_readdatavalid -> niosGe:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;       // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;    // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;          // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;           // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_niosge_debug_mem_slave_readdata;       // niosGe:debug_mem_slave_readdata -> mm_interconnect_0:niosGe_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosge_debug_mem_slave_waitrequest;    // niosGe:debug_mem_slave_waitrequest -> mm_interconnect_0:niosGe_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosge_debug_mem_slave_debugaccess;    // mm_interconnect_0:niosGe_debug_mem_slave_debugaccess -> niosGe:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosge_debug_mem_slave_address;        // mm_interconnect_0:niosGe_debug_mem_slave_address -> niosGe:debug_mem_slave_address
	wire         mm_interconnect_0_niosge_debug_mem_slave_read;           // mm_interconnect_0:niosGe_debug_mem_slave_read -> niosGe:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosge_debug_mem_slave_byteenable;     // mm_interconnect_0:niosGe_debug_mem_slave_byteenable -> niosGe:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosge_debug_mem_slave_write;          // mm_interconnect_0:niosGe_debug_mem_slave_write -> niosGe:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosge_debug_mem_slave_writedata;      // mm_interconnect_0:niosGe_debug_mem_slave_writedata -> niosGe:debug_mem_slave_writedata
	wire         mm_interconnect_0_flash_epcs_control_port_chipselect;    // mm_interconnect_0:flash_epcs_control_port_chipselect -> flash:chipselect
	wire  [31:0] mm_interconnect_0_flash_epcs_control_port_readdata;      // flash:readdata -> mm_interconnect_0:flash_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_flash_epcs_control_port_address;       // mm_interconnect_0:flash_epcs_control_port_address -> flash:address
	wire         mm_interconnect_0_flash_epcs_control_port_read;          // mm_interconnect_0:flash_epcs_control_port_read -> flash:read_n
	wire         mm_interconnect_0_flash_epcs_control_port_write;         // mm_interconnect_0:flash_epcs_control_port_write -> flash:write_n
	wire  [31:0] mm_interconnect_0_flash_epcs_control_port_writedata;     // mm_interconnect_0:flash_epcs_control_port_writedata -> flash:writedata
	wire         mm_interconnect_0_bl_n_s1_chipselect;                    // mm_interconnect_0:bl_n_s1_chipselect -> bl_n:chipselect
	wire  [31:0] mm_interconnect_0_bl_n_s1_readdata;                      // bl_n:readdata -> mm_interconnect_0:bl_n_s1_readdata
	wire   [1:0] mm_interconnect_0_bl_n_s1_address;                       // mm_interconnect_0:bl_n_s1_address -> bl_n:address
	wire         mm_interconnect_0_bl_n_s1_write;                         // mm_interconnect_0:bl_n_s1_write -> bl_n:write_n
	wire  [31:0] mm_interconnect_0_bl_n_s1_writedata;                     // mm_interconnect_0:bl_n_s1_writedata -> bl_n:writedata
	wire         mm_interconnect_0_bl_p_s1_chipselect;                    // mm_interconnect_0:bl_p_s1_chipselect -> bl_p:chipselect
	wire  [31:0] mm_interconnect_0_bl_p_s1_readdata;                      // bl_p:readdata -> mm_interconnect_0:bl_p_s1_readdata
	wire   [1:0] mm_interconnect_0_bl_p_s1_address;                       // mm_interconnect_0:bl_p_s1_address -> bl_p:address
	wire         mm_interconnect_0_bl_p_s1_write;                         // mm_interconnect_0:bl_p_s1_write -> bl_p:write_n
	wire  [31:0] mm_interconnect_0_bl_p_s1_writedata;                     // mm_interconnect_0:bl_p_s1_writedata -> bl_p:writedata
	wire         mm_interconnect_0_lcd_rd_s1_chipselect;                  // mm_interconnect_0:lcd_rd_s1_chipselect -> lcd_rd:chipselect
	wire  [31:0] mm_interconnect_0_lcd_rd_s1_readdata;                    // lcd_rd:readdata -> mm_interconnect_0:lcd_rd_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_rd_s1_address;                     // mm_interconnect_0:lcd_rd_s1_address -> lcd_rd:address
	wire         mm_interconnect_0_lcd_rd_s1_write;                       // mm_interconnect_0:lcd_rd_s1_write -> lcd_rd:write_n
	wire  [31:0] mm_interconnect_0_lcd_rd_s1_writedata;                   // mm_interconnect_0:lcd_rd_s1_writedata -> lcd_rd:writedata
	wire         mm_interconnect_0_lcd32_data_s1_chipselect;              // mm_interconnect_0:lcd32_data_s1_chipselect -> lcd32_data:chipselect
	wire  [31:0] mm_interconnect_0_lcd32_data_s1_readdata;                // lcd32_data:readdata -> mm_interconnect_0:lcd32_data_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd32_data_s1_address;                 // mm_interconnect_0:lcd32_data_s1_address -> lcd32_data:address
	wire         mm_interconnect_0_lcd32_data_s1_write;                   // mm_interconnect_0:lcd32_data_s1_write -> lcd32_data:write_n
	wire  [31:0] mm_interconnect_0_lcd32_data_s1_writedata;               // mm_interconnect_0:lcd32_data_s1_writedata -> lcd32_data:writedata
	wire         mm_interconnect_0_lcd_wr_s1_chipselect;                  // mm_interconnect_0:lcd_wr_s1_chipselect -> lcd_wr:chipselect
	wire  [31:0] mm_interconnect_0_lcd_wr_s1_readdata;                    // lcd_wr:readdata -> mm_interconnect_0:lcd_wr_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_wr_s1_address;                     // mm_interconnect_0:lcd_wr_s1_address -> lcd_wr:address
	wire         mm_interconnect_0_lcd_wr_s1_write;                       // mm_interconnect_0:lcd_wr_s1_write -> lcd_wr:write_n
	wire  [31:0] mm_interconnect_0_lcd_wr_s1_writedata;                   // mm_interconnect_0:lcd_wr_s1_writedata -> lcd_wr:writedata
	wire         mm_interconnect_0_reset_s1_chipselect;                   // mm_interconnect_0:reset_s1_chipselect -> reset:chipselect
	wire  [31:0] mm_interconnect_0_reset_s1_readdata;                     // reset:readdata -> mm_interconnect_0:reset_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_s1_address;                      // mm_interconnect_0:reset_s1_address -> reset:address
	wire         mm_interconnect_0_reset_s1_write;                        // mm_interconnect_0:reset_s1_write -> reset:write_n
	wire  [31:0] mm_interconnect_0_reset_s1_writedata;                    // mm_interconnect_0:reset_s1_writedata -> reset:writedata
	wire  [31:0] mm_interconnect_0_touch_irq_s1_readdata;                 // touch_irq:readdata -> mm_interconnect_0:touch_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_irq_s1_address;                  // mm_interconnect_0:touch_irq_s1_address -> touch_irq:address
	wire         mm_interconnect_0_lcd_rs_s1_chipselect;                  // mm_interconnect_0:lcd_rs_s1_chipselect -> lcd_rs:chipselect
	wire  [31:0] mm_interconnect_0_lcd_rs_s1_readdata;                    // lcd_rs:readdata -> mm_interconnect_0:lcd_rs_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_rs_s1_address;                     // mm_interconnect_0:lcd_rs_s1_address -> lcd_rs:address
	wire         mm_interconnect_0_lcd_rs_s1_write;                       // mm_interconnect_0:lcd_rs_s1_write -> lcd_rs:write_n
	wire  [31:0] mm_interconnect_0_lcd_rs_s1_writedata;                   // mm_interconnect_0:lcd_rs_s1_writedata -> lcd_rs:writedata
	wire         mm_interconnect_0_touch_cs_s1_chipselect;                // mm_interconnect_0:touch_cs_s1_chipselect -> touch_cs:chipselect
	wire  [31:0] mm_interconnect_0_touch_cs_s1_readdata;                  // touch_cs:readdata -> mm_interconnect_0:touch_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_cs_s1_address;                   // mm_interconnect_0:touch_cs_s1_address -> touch_cs:address
	wire         mm_interconnect_0_touch_cs_s1_write;                     // mm_interconnect_0:touch_cs_s1_write -> touch_cs:write_n
	wire  [31:0] mm_interconnect_0_touch_cs_s1_writedata;                 // mm_interconnect_0:touch_cs_s1_writedata -> touch_cs:writedata
	wire         mm_interconnect_0_lcd_cs_s1_chipselect;                  // mm_interconnect_0:lcd_cs_s1_chipselect -> lcd_cs:chipselect
	wire  [31:0] mm_interconnect_0_lcd_cs_s1_readdata;                    // lcd_cs:readdata -> mm_interconnect_0:lcd_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_cs_s1_address;                     // mm_interconnect_0:lcd_cs_s1_address -> lcd_cs:address
	wire         mm_interconnect_0_lcd_cs_s1_write;                       // mm_interconnect_0:lcd_cs_s1_write -> lcd_cs:write_n
	wire  [31:0] mm_interconnect_0_lcd_cs_s1_writedata;                   // mm_interconnect_0:lcd_cs_s1_writedata -> lcd_cs:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                   // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                     // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                      // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                        // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                    // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                        // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                         // mm_interconnect_0:SW_s1_address -> SW:address
	wire         mm_interconnect_0_led_s1_chipselect;                     // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                       // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                        // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_write;                          // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                      // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                   // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                     // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                  // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                      // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                         // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                   // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                        // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                    // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_spi_touch_spi_control_port_chipselect; // mm_interconnect_0:spi_touch_spi_control_port_chipselect -> spi_touch:spi_select
	wire  [15:0] mm_interconnect_0_spi_touch_spi_control_port_readdata;   // spi_touch:data_to_cpu -> mm_interconnect_0:spi_touch_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_touch_spi_control_port_address;    // mm_interconnect_0:spi_touch_spi_control_port_address -> spi_touch:mem_addr
	wire         mm_interconnect_0_spi_touch_spi_control_port_read;       // mm_interconnect_0:spi_touch_spi_control_port_read -> spi_touch:read_n
	wire         mm_interconnect_0_spi_touch_spi_control_port_write;      // mm_interconnect_0:spi_touch_spi_control_port_write -> spi_touch:write_n
	wire  [15:0] mm_interconnect_0_spi_touch_spi_control_port_writedata;  // mm_interconnect_0:spi_touch_spi_control_port_writedata -> spi_touch:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                // spi_touch:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver3_irq;                                // flash:irq -> irq_mapper:receiver3_irq
	wire  [31:0] niosge_irq_irq;                                          // irq_mapper:sender_irq -> niosGe:irq
	wire         irq_mapper_receiver1_irq;                                // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                           // jtag:av_irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                       // timer:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [LED:reset_n, SW:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, jtag:rst_n, mm_interconnect_0:jtag_reset_reset_bridge_in_reset_reset, timer:reset_n]
	wire         niosge_debug_reset_request_reset;                        // niosGe:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                      // rst_controller_001:reset_out -> [bl_n:reset_n, bl_p:reset_n, flash:reset_n, lcd32_data:reset_n, lcd_cs:reset_n, lcd_rd:reset_n, lcd_rs:reset_n, lcd_wr:reset_n, mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, reset:reset_n, rst_translator:in_reset, sysid:reset_n, touch_cs:reset_n, touch_irq:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                  // rst_controller_001:reset_req -> [flash:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                      // rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:niosGe_reset_reset_bridge_in_reset_reset, niosGe:reset_n, rst_translator_001:in_reset, sdram:reset_n, spi_touch:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                  // rst_controller_002:reset_req -> [niosGe:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                      // rst_controller_003:reset_out -> pll:reset

	mi_nios_LED led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	mi_nios_SW sw (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_export)                         // external_connection.export
	);

	mi_nios_bl_n bl_n (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_bl_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bl_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bl_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bl_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bl_n_s1_readdata),   //                    .readdata
		.out_port   (bl_n_export)                           // external_connection.export
	);

	mi_nios_bl_n bl_p (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_bl_p_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bl_p_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bl_p_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bl_p_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bl_p_s1_readdata),   //                    .readdata
		.out_port   (bl_p_export)                           // external_connection.export
	);

	mi_nios_flash flash (
		.clk        (pll_c0_clk),                                           //               clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //             reset.reset_n
		.reset_req  (rst_controller_001_reset_out_reset_req),               //                  .reset_req
		.address    (mm_interconnect_0_flash_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_flash_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_flash_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_flash_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_flash_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_flash_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver3_irq),                             //               irq.irq
		.dclk       (flash_dclk),                                           //          external.export
		.sce        (flash_sce),                                            //                  .export
		.sdo        (flash_sdo),                                            //                  .export
		.data0      (flash_data0)                                           //                  .export
	);

	mi_nios_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_receiver_irq)                         //               irq.irq
	);

	mi_nios_lcd32_data lcd32_data (
		.clk        (pll_c0_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lcd32_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd32_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd32_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd32_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd32_data_s1_readdata),   //                    .readdata
		.bidir_port (lcd32_data_export)                           // external_connection.export
	);

	mi_nios_bl_n lcd_cs (
		.clk        (pll_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_lcd_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_cs_s1_readdata),   //                    .readdata
		.out_port   (lcd_cs_export)                           // external_connection.export
	);

	mi_nios_bl_n lcd_rd (
		.clk        (pll_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_lcd_rd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_rd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_rd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_rd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_rd_s1_readdata),   //                    .readdata
		.out_port   (lcd_rd_export)                           // external_connection.export
	);

	mi_nios_bl_n lcd_rs (
		.clk        (pll_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_lcd_rs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_rs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_rs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_rs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_rs_s1_readdata),   //                    .readdata
		.out_port   (lcd_rs_export)                           // external_connection.export
	);

	mi_nios_bl_n lcd_wr (
		.clk        (pll_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_lcd_wr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_wr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_wr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_wr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_wr_s1_readdata),   //                    .readdata
		.out_port   (lcd_wr_export)                           // external_connection.export
	);

	mi_nios_niosGe niosge (
		.clk                                 (pll_c0_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                  //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),               //                          .reset_req
		.d_address                           (niosge_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosge_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosge_data_master_read),                              //                          .read
		.d_readdata                          (niosge_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosge_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosge_data_master_write),                             //                          .write
		.d_writedata                         (niosge_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (niosge_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (niosge_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosge_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosge_instruction_master_read),                       //                          .read
		.i_readdata                          (niosge_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosge_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (niosge_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (niosge_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (niosge_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosge_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosge_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosge_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosge_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosge_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosge_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosge_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosge_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	mi_nios_pll pll (
		.clk       (clk_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_003_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (pll_c0_clk),                         //                    c0.clk
		.c1        (sdram_clk_clk),                      //                    c1.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	mi_nios_bl_n reset (
		.clk        (pll_c0_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_s1_readdata),   //                    .readdata
		.out_port   (reset_1_export)                         // external_connection.export
	);

	mi_nios_sdram sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	mi_nios_spi_touch spi_touch (
		.clk           (pll_c0_clk),                                              //              clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_touch_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_touch_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_touch_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_touch_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_touch_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_touch_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver0_irq),                                //              irq.irq
		.MISO          (spi_touch_MISO),                                          //         external.export
		.MOSI          (spi_touch_MOSI),                                          //                 .export
		.SCLK          (spi_touch_SCLK),                                          //                 .export
		.SS_n          (spi_touch_SS_n)                                           //                 .export
	);

	mi_nios_sysid sysid (
		.clock    (pll_c0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	mi_nios_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)      //   irq.irq
	);

	mi_nios_bl_n touch_cs (
		.clk        (pll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_touch_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_cs_s1_readdata),   //                    .readdata
		.out_port   (touch_cs_export)                           // external_connection.export
	);

	mi_nios_touch_irq touch_irq (
		.clk      (pll_c0_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_touch_irq_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_touch_irq_s1_readdata), //                    .readdata
		.in_port  (touch_irq_export)                         // external_connection.export
	);

	mi_nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                           (clk_clk),                                                 //                         clk_50_clk.clk
		.pll_c0_clk                               (pll_c0_clk),                                              //                             pll_c0.clk
		.jtag_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                          //   jtag_reset_reset_bridge_in_reset.reset
		.niosGe_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                      // niosGe_reset_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                      //  sysid_reset_reset_bridge_in_reset.reset
		.niosGe_data_master_address               (niosge_data_master_address),                              //                 niosGe_data_master.address
		.niosGe_data_master_waitrequest           (niosge_data_master_waitrequest),                          //                                   .waitrequest
		.niosGe_data_master_byteenable            (niosge_data_master_byteenable),                           //                                   .byteenable
		.niosGe_data_master_read                  (niosge_data_master_read),                                 //                                   .read
		.niosGe_data_master_readdata              (niosge_data_master_readdata),                             //                                   .readdata
		.niosGe_data_master_readdatavalid         (niosge_data_master_readdatavalid),                        //                                   .readdatavalid
		.niosGe_data_master_write                 (niosge_data_master_write),                                //                                   .write
		.niosGe_data_master_writedata             (niosge_data_master_writedata),                            //                                   .writedata
		.niosGe_data_master_debugaccess           (niosge_data_master_debugaccess),                          //                                   .debugaccess
		.niosGe_instruction_master_address        (niosge_instruction_master_address),                       //          niosGe_instruction_master.address
		.niosGe_instruction_master_waitrequest    (niosge_instruction_master_waitrequest),                   //                                   .waitrequest
		.niosGe_instruction_master_read           (niosge_instruction_master_read),                          //                                   .read
		.niosGe_instruction_master_readdata       (niosge_instruction_master_readdata),                      //                                   .readdata
		.niosGe_instruction_master_readdatavalid  (niosge_instruction_master_readdatavalid),                 //                                   .readdatavalid
		.bl_n_s1_address                          (mm_interconnect_0_bl_n_s1_address),                       //                            bl_n_s1.address
		.bl_n_s1_write                            (mm_interconnect_0_bl_n_s1_write),                         //                                   .write
		.bl_n_s1_readdata                         (mm_interconnect_0_bl_n_s1_readdata),                      //                                   .readdata
		.bl_n_s1_writedata                        (mm_interconnect_0_bl_n_s1_writedata),                     //                                   .writedata
		.bl_n_s1_chipselect                       (mm_interconnect_0_bl_n_s1_chipselect),                    //                                   .chipselect
		.bl_p_s1_address                          (mm_interconnect_0_bl_p_s1_address),                       //                            bl_p_s1.address
		.bl_p_s1_write                            (mm_interconnect_0_bl_p_s1_write),                         //                                   .write
		.bl_p_s1_readdata                         (mm_interconnect_0_bl_p_s1_readdata),                      //                                   .readdata
		.bl_p_s1_writedata                        (mm_interconnect_0_bl_p_s1_writedata),                     //                                   .writedata
		.bl_p_s1_chipselect                       (mm_interconnect_0_bl_p_s1_chipselect),                    //                                   .chipselect
		.flash_epcs_control_port_address          (mm_interconnect_0_flash_epcs_control_port_address),       //            flash_epcs_control_port.address
		.flash_epcs_control_port_write            (mm_interconnect_0_flash_epcs_control_port_write),         //                                   .write
		.flash_epcs_control_port_read             (mm_interconnect_0_flash_epcs_control_port_read),          //                                   .read
		.flash_epcs_control_port_readdata         (mm_interconnect_0_flash_epcs_control_port_readdata),      //                                   .readdata
		.flash_epcs_control_port_writedata        (mm_interconnect_0_flash_epcs_control_port_writedata),     //                                   .writedata
		.flash_epcs_control_port_chipselect       (mm_interconnect_0_flash_epcs_control_port_chipselect),    //                                   .chipselect
		.jtag_avalon_jtag_slave_address           (mm_interconnect_0_jtag_avalon_jtag_slave_address),        //             jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write             (mm_interconnect_0_jtag_avalon_jtag_slave_write),          //                                   .write
		.jtag_avalon_jtag_slave_read              (mm_interconnect_0_jtag_avalon_jtag_slave_read),           //                                   .read
		.jtag_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),       //                                   .readdata
		.jtag_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),      //                                   .writedata
		.jtag_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),    //                                   .waitrequest
		.jtag_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),     //                                   .chipselect
		.lcd32_data_s1_address                    (mm_interconnect_0_lcd32_data_s1_address),                 //                      lcd32_data_s1.address
		.lcd32_data_s1_write                      (mm_interconnect_0_lcd32_data_s1_write),                   //                                   .write
		.lcd32_data_s1_readdata                   (mm_interconnect_0_lcd32_data_s1_readdata),                //                                   .readdata
		.lcd32_data_s1_writedata                  (mm_interconnect_0_lcd32_data_s1_writedata),               //                                   .writedata
		.lcd32_data_s1_chipselect                 (mm_interconnect_0_lcd32_data_s1_chipselect),              //                                   .chipselect
		.lcd_cs_s1_address                        (mm_interconnect_0_lcd_cs_s1_address),                     //                          lcd_cs_s1.address
		.lcd_cs_s1_write                          (mm_interconnect_0_lcd_cs_s1_write),                       //                                   .write
		.lcd_cs_s1_readdata                       (mm_interconnect_0_lcd_cs_s1_readdata),                    //                                   .readdata
		.lcd_cs_s1_writedata                      (mm_interconnect_0_lcd_cs_s1_writedata),                   //                                   .writedata
		.lcd_cs_s1_chipselect                     (mm_interconnect_0_lcd_cs_s1_chipselect),                  //                                   .chipselect
		.lcd_rd_s1_address                        (mm_interconnect_0_lcd_rd_s1_address),                     //                          lcd_rd_s1.address
		.lcd_rd_s1_write                          (mm_interconnect_0_lcd_rd_s1_write),                       //                                   .write
		.lcd_rd_s1_readdata                       (mm_interconnect_0_lcd_rd_s1_readdata),                    //                                   .readdata
		.lcd_rd_s1_writedata                      (mm_interconnect_0_lcd_rd_s1_writedata),                   //                                   .writedata
		.lcd_rd_s1_chipselect                     (mm_interconnect_0_lcd_rd_s1_chipselect),                  //                                   .chipselect
		.lcd_rs_s1_address                        (mm_interconnect_0_lcd_rs_s1_address),                     //                          lcd_rs_s1.address
		.lcd_rs_s1_write                          (mm_interconnect_0_lcd_rs_s1_write),                       //                                   .write
		.lcd_rs_s1_readdata                       (mm_interconnect_0_lcd_rs_s1_readdata),                    //                                   .readdata
		.lcd_rs_s1_writedata                      (mm_interconnect_0_lcd_rs_s1_writedata),                   //                                   .writedata
		.lcd_rs_s1_chipselect                     (mm_interconnect_0_lcd_rs_s1_chipselect),                  //                                   .chipselect
		.lcd_wr_s1_address                        (mm_interconnect_0_lcd_wr_s1_address),                     //                          lcd_wr_s1.address
		.lcd_wr_s1_write                          (mm_interconnect_0_lcd_wr_s1_write),                       //                                   .write
		.lcd_wr_s1_readdata                       (mm_interconnect_0_lcd_wr_s1_readdata),                    //                                   .readdata
		.lcd_wr_s1_writedata                      (mm_interconnect_0_lcd_wr_s1_writedata),                   //                                   .writedata
		.lcd_wr_s1_chipselect                     (mm_interconnect_0_lcd_wr_s1_chipselect),                  //                                   .chipselect
		.LED_s1_address                           (mm_interconnect_0_led_s1_address),                        //                             LED_s1.address
		.LED_s1_write                             (mm_interconnect_0_led_s1_write),                          //                                   .write
		.LED_s1_readdata                          (mm_interconnect_0_led_s1_readdata),                       //                                   .readdata
		.LED_s1_writedata                         (mm_interconnect_0_led_s1_writedata),                      //                                   .writedata
		.LED_s1_chipselect                        (mm_interconnect_0_led_s1_chipselect),                     //                                   .chipselect
		.niosGe_debug_mem_slave_address           (mm_interconnect_0_niosge_debug_mem_slave_address),        //             niosGe_debug_mem_slave.address
		.niosGe_debug_mem_slave_write             (mm_interconnect_0_niosge_debug_mem_slave_write),          //                                   .write
		.niosGe_debug_mem_slave_read              (mm_interconnect_0_niosge_debug_mem_slave_read),           //                                   .read
		.niosGe_debug_mem_slave_readdata          (mm_interconnect_0_niosge_debug_mem_slave_readdata),       //                                   .readdata
		.niosGe_debug_mem_slave_writedata         (mm_interconnect_0_niosge_debug_mem_slave_writedata),      //                                   .writedata
		.niosGe_debug_mem_slave_byteenable        (mm_interconnect_0_niosge_debug_mem_slave_byteenable),     //                                   .byteenable
		.niosGe_debug_mem_slave_waitrequest       (mm_interconnect_0_niosge_debug_mem_slave_waitrequest),    //                                   .waitrequest
		.niosGe_debug_mem_slave_debugaccess       (mm_interconnect_0_niosge_debug_mem_slave_debugaccess),    //                                   .debugaccess
		.reset_s1_address                         (mm_interconnect_0_reset_s1_address),                      //                           reset_s1.address
		.reset_s1_write                           (mm_interconnect_0_reset_s1_write),                        //                                   .write
		.reset_s1_readdata                        (mm_interconnect_0_reset_s1_readdata),                     //                                   .readdata
		.reset_s1_writedata                       (mm_interconnect_0_reset_s1_writedata),                    //                                   .writedata
		.reset_s1_chipselect                      (mm_interconnect_0_reset_s1_chipselect),                   //                                   .chipselect
		.sdram_s1_address                         (mm_interconnect_0_sdram_s1_address),                      //                           sdram_s1.address
		.sdram_s1_write                           (mm_interconnect_0_sdram_s1_write),                        //                                   .write
		.sdram_s1_read                            (mm_interconnect_0_sdram_s1_read),                         //                                   .read
		.sdram_s1_readdata                        (mm_interconnect_0_sdram_s1_readdata),                     //                                   .readdata
		.sdram_s1_writedata                       (mm_interconnect_0_sdram_s1_writedata),                    //                                   .writedata
		.sdram_s1_byteenable                      (mm_interconnect_0_sdram_s1_byteenable),                   //                                   .byteenable
		.sdram_s1_readdatavalid                   (mm_interconnect_0_sdram_s1_readdatavalid),                //                                   .readdatavalid
		.sdram_s1_waitrequest                     (mm_interconnect_0_sdram_s1_waitrequest),                  //                                   .waitrequest
		.sdram_s1_chipselect                      (mm_interconnect_0_sdram_s1_chipselect),                   //                                   .chipselect
		.spi_touch_spi_control_port_address       (mm_interconnect_0_spi_touch_spi_control_port_address),    //         spi_touch_spi_control_port.address
		.spi_touch_spi_control_port_write         (mm_interconnect_0_spi_touch_spi_control_port_write),      //                                   .write
		.spi_touch_spi_control_port_read          (mm_interconnect_0_spi_touch_spi_control_port_read),       //                                   .read
		.spi_touch_spi_control_port_readdata      (mm_interconnect_0_spi_touch_spi_control_port_readdata),   //                                   .readdata
		.spi_touch_spi_control_port_writedata     (mm_interconnect_0_spi_touch_spi_control_port_writedata),  //                                   .writedata
		.spi_touch_spi_control_port_chipselect    (mm_interconnect_0_spi_touch_spi_control_port_chipselect), //                                   .chipselect
		.SW_s1_address                            (mm_interconnect_0_sw_s1_address),                         //                              SW_s1.address
		.SW_s1_readdata                           (mm_interconnect_0_sw_s1_readdata),                        //                                   .readdata
		.sysid_control_slave_address              (mm_interconnect_0_sysid_control_slave_address),           //                sysid_control_slave.address
		.sysid_control_slave_readdata             (mm_interconnect_0_sysid_control_slave_readdata),          //                                   .readdata
		.timer_s1_address                         (mm_interconnect_0_timer_s1_address),                      //                           timer_s1.address
		.timer_s1_write                           (mm_interconnect_0_timer_s1_write),                        //                                   .write
		.timer_s1_readdata                        (mm_interconnect_0_timer_s1_readdata),                     //                                   .readdata
		.timer_s1_writedata                       (mm_interconnect_0_timer_s1_writedata),                    //                                   .writedata
		.timer_s1_chipselect                      (mm_interconnect_0_timer_s1_chipselect),                   //                                   .chipselect
		.touch_cs_s1_address                      (mm_interconnect_0_touch_cs_s1_address),                   //                        touch_cs_s1.address
		.touch_cs_s1_write                        (mm_interconnect_0_touch_cs_s1_write),                     //                                   .write
		.touch_cs_s1_readdata                     (mm_interconnect_0_touch_cs_s1_readdata),                  //                                   .readdata
		.touch_cs_s1_writedata                    (mm_interconnect_0_touch_cs_s1_writedata),                 //                                   .writedata
		.touch_cs_s1_chipselect                   (mm_interconnect_0_touch_cs_s1_chipselect),                //                                   .chipselect
		.touch_irq_s1_address                     (mm_interconnect_0_touch_irq_s1_address),                  //                       touch_irq_s1.address
		.touch_irq_s1_readdata                    (mm_interconnect_0_touch_irq_s1_readdata)                  //                                   .readdata
	);

	mi_nios_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (niosge_irq_irq)                      //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                   // reset_in0.reset
		.reset_in1      (niosge_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (niosge_debug_reset_request_reset),       // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
